library verilog;
use verilog.vl_types.all;
entity lab06_all_vlg_tst is
end lab06_all_vlg_tst;
