library verilog;
use verilog.vl_types.all;
entity ID_EX is
    port(
        clk             : in     vl_logic;
        PC_src          : in     vl_logic_vector(1 downto 0);
        Regwr           : in     vl_logic;
        regdst          : in     vl_logic_vector(1 downto 0);
        MemOp           : in     vl_logic_vector(2 downto 0);
        CacheOp         : in     vl_logic_vector(2 downto 0);
        Choice          : in     vl_logic;
        Rd              : in     vl_logic_vector(4 downto 0);
        Rs              : in     vl_logic_vector(4 downto 0);
        Rt              : in     vl_logic_vector(4 downto 0);
        Mem_byte_wr_in  : in     vl_logic_vector(3 downto 0);
        MemRead         : in     vl_logic;
        Extend          : in     vl_logic_vector(1 downto 0);
        branch          : in     vl_logic;
        Jump            : in     vl_logic;
        Condition       : in     vl_logic_vector(2 downto 0);
        ExResultSrc     : in     vl_logic_vector(2 downto 0);
        ALUSrcA         : in     vl_logic;
        ALUSrcB         : in     vl_logic;
        ALU_op          : in     vl_logic_vector(3 downto 0);
        Shift_amountSrc : in     vl_logic;
        Shift_op        : in     vl_logic_vector(1 downto 0);
        Immediate32     : in     vl_logic_vector(31 downto 0);
        OperandA        : in     vl_logic_vector(31 downto 0);
        OperandB        : in     vl_logic_vector(31 downto 0);
        WBtype          : in     vl_logic_vector(3 downto 0);
        add_pc          : in     vl_logic_vector(31 downto 0);
        Regwr2          : out    vl_logic;
        regdst2         : out    vl_logic_vector(1 downto 0);
        MemOp2          : out    vl_logic_vector(2 downto 0);
        CacheOp2        : out    vl_logic_vector(2 downto 0);
        Choice2         : out    vl_logic;
        Rd2             : out    vl_logic_vector(4 downto 0);
        Rs2             : out    vl_logic_vector(4 downto 0);
        Rt2             : out    vl_logic_vector(4 downto 0);
        Mem_byte_wr_in2 : out    vl_logic_vector(3 downto 0);
        MemRead2        : out    vl_logic;
        Extend2         : out    vl_logic_vector(1 downto 0);
        branch2         : out    vl_logic;
        Jump2           : out    vl_logic;
        Condition2      : out    vl_logic_vector(2 downto 0);
        ExResultSrc2    : out    vl_logic_vector(2 downto 0);
        ALUSrcA2        : out    vl_logic;
        ALUSrcB2        : out    vl_logic;
        ALU_op2         : out    vl_logic_vector(3 downto 0);
        Shift_amountSrc2: out    vl_logic;
        Shift_op2       : out    vl_logic_vector(1 downto 0);
        Immediate32_2   : out    vl_logic_vector(31 downto 0);
        OperandA2       : out    vl_logic_vector(31 downto 0);
        OperandB2       : out    vl_logic_vector(31 downto 0);
        WBtype2         : out    vl_logic_vector(3 downto 0);
        add_pc2         : out    vl_logic_vector(31 downto 0)
    );
end ID_EX;
